module alsu_tb();

reg [2:0] A, B, opcode;
reg cin,
      serial_in,
      direction,
      red_op_A,
      red_op_B,
      bypass_A,
      bypass_B,
      clk,
      rst;
wire [5:0] out;
wire [15:0] leds;



endmodule