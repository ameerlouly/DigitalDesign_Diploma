module Q3_adder(A, B, C);

    input [3:0] A, B;
    output [3:0] C;

    assign C = A + B;

endmodule