module alu(A, B,  opcode, rst, clk, out);


endmodule