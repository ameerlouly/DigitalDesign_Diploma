module simple_dsp();

endmodule